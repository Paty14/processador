library verilog;
use verilog.vl_types.all;
entity testeIntegracao is
end testeIntegracao;
