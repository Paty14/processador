library verilog;
use verilog.vl_types.all;
entity zzzTesteMemoria is
end zzzTesteMemoria;
